module testElement(out, in);
input in;
output out;

wire   w;

assign w = in;
assign out = w;

endmodule
